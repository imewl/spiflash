//---------------------------------------------------------------------
//                                          
//     ____     ____     _____    _____    __  __    _____     ____  
//    /\___\   /\___\   /\____\  |\_____\ |\_\|\_\  |\____\   /\___\ 
//   |\/ _ _\ |\/ _  \  \/ ____| ||  ___| ||  \/  | \|_   _| |\/ _ _\
//   || |     || /_\  | \| |__   || |_\   ||      |   || |   || |    
//   || |___  || |__| |  _\__ \  ||  _|_  || |\/| |  _|| |_  || |___ 
//   \| |___\ || | || | |\__\| | || |___\ || |  | | |\_| |_\ \| |___\
//    \\____/ \|_| \|_| \|____/  \|_____| \|_|  |_| \|_____|  \\____/
//
//  COPYRIGHT 2017, ALL RIGHTS RESERVED
//  
//  Filename:   qspi_controller
//  Author:          
//  Date:            
//
//  Project:         
//  Descriptions: AHB Interface register for Quad-SPI controller.
//---------------------------------------------------------------------
module qspi_controller (
                // AHB Slave Interface
				ahb_rst_i,
                ahb_clk_i,
				
						);
//--------------------------------
//  Ports
//--------------------------------
input           ahb_rst_i;
input           ahb_clk_i;


//--------------------------------
//  Wires and REGs
//--------------------------------

endmodule
